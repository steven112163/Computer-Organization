`timescale 1ns / 1ps
//Subject:     CO project 3 - Adder
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      0510002 �K౳� 0510009 �i౸�
//--------------------------------------------------------------------------------
//Date:        2018/05/11
//--------------------------------------------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Adder(
    src1_i,  //32 bit src1_i (input)
	src2_i,  //32 bit src2_i (input)
	sum_o    //32 bit sum_o  (output)
	);
     
//I/O ports
input   [31:0] src1_i;
input   [31:0] src2_i;
output  [31:0] sum_o;

//Internal Signals
reg     [31:0] sum_o;

//Main function
always@ (*) begin
	sum_o <= src1_i + src2_i;
end

endmodule